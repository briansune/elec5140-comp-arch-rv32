`define N_EXT_INTS 24

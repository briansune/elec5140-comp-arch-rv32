parameter risc_v2udp_ack	= {"a","c","k","+"};
parameter risc_v2udp_OK		= {"O","K","!","\n"};
parameter risc_v2udp_ERROR	= {"E","R","!","\n"};

parameter udp2risc_v_nop	= {"n","o","p","-"};
parameter udp2risc_v_rst	= {"r","s","t","-"};
parameter udp2risc_v_prg	= {"p","r","g","-"};
parameter udp2risc_v_run	= {"r","u","n","-"};
parameter udp2risc_v_held	= {"h","l","d","-"};
parameter udp2risc_v_RROM	= {"r","d","\0","\0"};





`define MEM_BUS_WIDTH  32
`define MEM_BUS_NBYTES  4
`define MEM_ADDR_WIDTH 32

`define MEM_TRANS_WIDTH 2
`define MEM_TRANS_IDLE   `MEM_TRANS_WIDTH'd0
`define MEM_TRANS_BUSY   `MEM_TRANS_WIDTH'd1
`define MEM_TRANS_NONSEQ `MEM_TRANS_WIDTH'd2
`define MEM_TRANS_SEQ    `MEM_TRANS_WIDTH'd3

`define MEM_PROT_WIDTH 4
`define MEM_NO_PROT `MEM_PROT_WIDTH'd0

`define MEM_BURST_WIDTH 3
`define MEM_BURST_SINGLE `MEM_BURST_WIDTH'd0

`define MEM_MASTER_NO_LOCK 1'b0

`define MEM_RESP_WIDTH 1
`define MEM_RESP_OKAY  `MEM_RESP_WIDTH'd0
`define MEM_RESP_ERROR `MEM_RESP_WIDTH'd1

`define MEM_SIZE_WIDTH 3
`define MEM_SIZE_BYTE     `MEM_SIZE_WIDTH'd0
`define MEM_SIZE_HALFWORD `MEM_SIZE_WIDTH'd1
`define MEM_SIZE_WORD     `MEM_SIZE_WIDTH'd2
